library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
USE ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use work.mes_composants.all;

entity genHL is
generic( N_div : natural := 250);
    Port ( clk : in STD_LOGIC;
           reset : in STD_LOGIC;
           enRead : out STD_LOGIC;
           enWrite : out  std_logic
           );
end genHL;

architecture genHl of genHL is
    signal cpt1:std_logic_vector(7 downto 0):=(others=>'0');
    signal impulsion,raz : STD_LOGIC := '0';
    
begin
  DCPT_M1 : DCPT_M generic map(8)
    port map (
            enable => '1',
            ud     => '0',
            clk    => clk,
            reset  => raz,
            cptr   => cpt1
        );
                   
  impulsion <='1' when cpt1 = CONV_STD_LOGIC_VECTOR(N_div,8) else '0';
  raz <='1' when reset='1' or impulsion='1' else '0';
  
  enRead<=impulsion;
  enWrite<=not impulsion;   
end;

